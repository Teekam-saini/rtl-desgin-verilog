//conflict branch: expermenting with and gate
module and_gate(a,b,c,y);

 input a,b,c;
 output y;

 assign y = a&b&c;

endmodule

